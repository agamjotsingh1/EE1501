module loop_adder (
);

endmodule
